library verilog;
use verilog.vl_types.all;
entity DES_Testbench is
end DES_Testbench;
